//`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////////
//// Company: 
//// Engineer: 
//// 
//// Create Date: 04.03.2024 01:38:33
//// Design Name: 
//// Module Name: decoder4x16_testbench
//// Project Name: 
//// Target Devices: 
//// Tool Versions: 
//// Description: 
//// 
//// Dependencies: 
//// 
//// Revision:
//// Revision 0.01 - File Created
//// Additional Comments:
//// 
////////////////////////////////////////////////////////////////////////////////////


//module decoder4x16_testbench();

//reg A, B, C, D;
//wire [15:0] O;

//decoder_4x16_enable dut(A,B,C,D,O);
//initial begin
//        {A,B,C,D} = 4'b0001;
//        #10
//        {A,B,C,D} = 4'b0011;
//        #10
//        {A,B,C,D} = 4'b1001;
//        #10
//        {A,B,C,D} = 4'b1111;
//        #10
        
//        $finish;
//        end
//endmodule